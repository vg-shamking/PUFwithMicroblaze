library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package parameters is

    constant C_LENGTH : natural :=32;
    constant C_DFF_TYPE : string := "PRIMITIVE";
    
    alias sl is STD_LOGIC ;
    alias slv is STD_LOGIC_VECTOR ;

end package;
